library ieee;
use ieee.std_logic_1164.all;

entity io is
end entity;

architecture one of io is
begin
end entity;